`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: University of Stuttgart, ITI
// Engineer: Alexander Kharitonov
// 
// Create Date: 29.06.2023 15:45:28
// Design Name: 
// Module Name: soc_registers
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: Defines for SoC peripheral registers.
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`ifndef SOC_REGISTERS_HEADER //include guard
`define SOC_REGISTERS_HEADER



//**************************** GENERAL ****************************
//Register access types
`define REG_TYPE_MAIN 2'd0
`define REG_TYPE_SET 2'd1
`define REG_TYPE_CLR 2'd2
`define REG_TYPE_INV 2'd3

//Register access type implementation macro
`define REG_WRITEVAL(current, write, type) (\
    (type == `REG_TYPE_MAIN) ? (write) : (\
    (type == `REG_TYPE_SET) ? ((current) | (write)) : (\
    (type == `REG_TYPE_CLR) ? ((current) & ~(write)) : (\
    ((current) ^ (write))))))



//**************************** SOC CONTROL ****************************
`define REG_SOCCTL_CONTROL      8'h00 //control register - core halt, core reset, soc reset, interrupt global en, control flags
`define REG_SOCCTL_INT_EN       8'h01 //enabled interrupts
`define REG_SOCCTL_INT_FLAGS    8'h02 //asserted interrupts



//**************************** GPIO ****************************
`define REG_GPIO_PORT           4'h0 //port register - pin status
`define REG_GPIO_LATCH          4'h1 //latch register - values outputted on output pins
`define REG_GPIO_DIR            4'h2 //direction register - pin directions (0 = input, 1 = output)
`define REG_GPIO_CNR            4'h3 //change notification enable - rising edge
`define REG_GPIO_CNF            4'h4 //change notification enable - falling edge
`define REG_GPIO_CN_STATE       4'h5 //change notification state - 1 if change occurred
`define REG_GPIO_INT_STATUS     4'hF //interrupt status - 1 if interrupt generated by given port



//**************************** PWM ****************************
`define REG_PWM_CONTROL         4'h0
`define REG_PWM_VALUE           4'h1
`define REG_PWM_NEXT_VALUE      4'h2



//**************************** TIMER ****************************
`define REG_TIMER_CONTROL       4'h0
`define REG_TIMER_COUNT         4'h1
`define REG_TIMER_PERIOD        4'h2
`define REG_TIMER_INT_STATUS    4'hF



`endif //include guard