----------------------------------------------------------------------------------
-- Company: Digilent
-- Engineer: Arthur Brown
-- 
--
-- Create Date:    13:01:51 02/15/2013 
-- Project Name:   pmodvga
-- Target Devices: arty
-- Tool versions:  2016.4
-- Additional Comments: 
--
-- Copyright Digilent 2017
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity vga_digilent is
    Port ( pxl_clk : in  STD_LOGIC;           
           VGA_HS_O : out  STD_LOGIC;
           VGA_VS_O : out  STD_LOGIC;
           PIXEL_I : in STD_LOGIC_VECTOR (7 downto 0);
           VGA_R : out  STD_LOGIC_VECTOR (3 downto 0);
           VGA_B : out  STD_LOGIC_VECTOR (3 downto 0);
           VGA_G : out  STD_LOGIC_VECTOR (3 downto 0);
           PXL_ADR_O : out STD_LOGIC_VECTOR (31 downto 0));
end vga_digilent;

architecture Behavioral of vga_digilent is

--Sync Generation constants

--***640x480@60Hz***--  Requires 25 MHz clock
constant FRAME_WIDTH : natural := 640;
constant FRAME_HEIGHT : natural := 480;
constant FRAME_H_START : natural := 60;

constant H_FP : natural := 16; --H front porch width (pixels)
constant H_PW : natural := 96; --H sync pulse width (pixels)
constant H_MAX : natural := 800; --H total period (pixels)

constant V_FP : natural := 10; --V front porch width (lines)
constant V_PW : natural := 2; --V sync pulse width (lines)
constant V_MAX : natural := 525; --V total period (lines)

--active <= '1' when h_cntr_reg >= 144 and h_cntr_reg <= 784 and v_cntr_reg >= 95 and v_cntr_reg <= 455 else
constant FIRST_COL : natural := 144; --First Horizontal Pixel in Frame
constant LAST_COL : natural := 784; --Last Horizontal Pixel in Frame
constant FIRST_LINE : natural := 95; --First line in Frame (+60px since we display 640x360)
constant LAST_LINE : natural := 455; --Last line in Frame (-60px since we display 640x360)

constant H_POL : std_logic := '0';
constant V_POL : std_logic := '0';

----***800x600@60Hz***--  Requires 40 MHz clock
--constant FRAME_WIDTH : natural := 800;
--constant FRAME_HEIGHT : natural := 600;
--
--constant H_FP : natural := 40; --H front porch width (pixels)
--constant H_PW : natural := 128; --H sync pulse width (pixels)
--constant H_MAX : natural := 1056; --H total period (pixels)
--
--constant V_FP : natural := 1; --V front porch width (lines)
--constant V_PW : natural := 4; --V sync pulse width (lines)
--constant V_MAX : natural := 628; --V total period (lines)
--
--constant H_POL : std_logic := '1';
--constant V_POL : std_logic := '1';


----***1280x720@60Hz***-- Requires 74.25 MHz clock
--constant FRAME_WIDTH : natural := 1280;
--constant FRAME_HEIGHT : natural := 720;
--
--constant H_FP : natural := 110; --H front porch width (pixels)
--constant H_PW : natural := 40; --H sync pulse width (pixels)
--constant H_MAX : natural := 1650; --H total period (pixels)
--
--constant V_FP : natural := 5; --V front porch width (lines)
--constant V_PW : natural := 5; --V sync pulse width (lines)
--constant V_MAX : natural := 750; --V total period (lines)
--
--constant H_POL : std_logic := '1';
--constant V_POL : std_logic := '1';

----***1280x1024@60Hz***-- Requires 108 MHz clock
--constant FRAME_WIDTH : natural := 1280;
--constant FRAME_HEIGHT : natural := 1024;

--constant H_FP : natural := 48; --H front porch width (pixels)
--constant H_PW : natural := 112; --H sync pulse width (pixels)
--constant H_MAX : natural := 1688; --H total period (pixels)

--constant V_FP : natural := 1; --V front porch width (lines)
--constant V_PW : natural := 3; --V sync pulse width (lines)
--constant V_MAX : natural := 1066; --V total period (lines)

--constant H_POL : std_logic := '1';
--constant V_POL : std_logic := '1';

----***1920x1080@60Hz***-- Requires 148.5 MHz pxl_clk
--constant FRAME_WIDTH : natural := 1920;
--constant FRAME_HEIGHT : natural := 1080;

--constant H_FP : natural := 88; --H front porch width (pixels)
--constant H_PW : natural := 44; --H sync pulse width (pixels)
--constant H_MAX : natural := 2200; --H total period (pixels)

--constant V_FP : natural := 4; --V front porch width (lines)
--constant V_PW : natural := 5; --V sync pulse width (lines)
--constant V_MAX : natural := 1125; --V total period (lines)

--constant H_POL : std_logic := '1';
--constant V_POL : std_logic := '1';

----Moving Box constants
--constant BOX_WIDTH : natural := 8;
--constant BOX_CLK_DIV : natural := 1000000; --MAX=(2^25 - 1)

--constant BOX_X_MAX : natural := (512 - BOX_WIDTH);
--constant BOX_Y_MAX : natural := (FRAME_HEIGHT - BOX_WIDTH);

--constant BOX_X_MIN : natural := 0;
--constant BOX_Y_MIN : natural := 256;

--constant BOX_X_INIT : std_logic_vector(11 downto 0) := x"000";
--constant BOX_Y_INIT : std_logic_vector(11 downto 0) := x"190"; --400

--signal pxl_clk : std_logic;
--signal active : std_logic;
signal active : std_logic := '0';

signal h_cntr_reg : std_logic_vector(11 downto 0) := (others =>'0');
signal v_cntr_reg : std_logic_vector(11 downto 0) := (others =>'0');
signal pxl_adr    : std_logic_vector(31 downto 0) := (others =>'0');
signal h_sync_reg : std_logic := not(H_POL);
signal v_sync_reg : std_logic := not(V_POL);

signal h_sync_dly_reg : std_logic := not(H_POL);
signal v_sync_dly_reg : std_logic :=  not(V_POL);

--signal vga_red_reg : std_logic_vector(3 downto 0) := (others =>'0');
--signal vga_green_reg : std_logic_vector(3 downto 0) := (others =>'0');
--signal vga_blue_reg : std_logic_vector(3 downto 0) := (others =>'0');

--signal vga_red : std_logic_vector(3 downto 0);
--signal vga_green : std_logic_vector(3 downto 0);
--signal vga_blue : std_logic_vector(3 downto 0);

--signal box_x_reg : std_logic_vector(11 downto 0) := BOX_X_INIT;
--signal box_x_dir : std_logic := '1';
--signal box_y_reg : std_logic_vector(11 downto 0) := BOX_Y_INIT;
--signal box_y_dir : std_logic := '1';
--signal box_cntr_reg : std_logic_vector(24 downto 0) := (others =>'0');

--signal update_box : std_logic;
--signal pixel_in_box : std_logic;


begin
  
   
--clk_div_inst : clk_wiz_0
--  port map
--   (-- Clock in ports
--    CLK_IN1 => CLK_I,
--    -- Clock out ports
--    CLK_OUT1 => pxl_clk);

  
  ----------------------------------------------------
  -------         TEST PATTERN LOGIC           -------
  ----------------------------------------------------
--  vga_red <= h_cntr_reg(5 downto 2) when (active = '1' and ((h_cntr_reg < 512 and v_cntr_reg < 256) and h_cntr_reg(8) = '1')) else
--              (others=>'1')         when (active = '1' and ((h_cntr_reg < 512 and not(v_cntr_reg < 256)) and not(pixel_in_box = '1'))) else
--              (others=>'1')         when (active = '1' and ((not(h_cntr_reg < 512) and (v_cntr_reg(8) = '1' and h_cntr_reg(3) = '1')) or
--                                          (not(h_cntr_reg < 512) and (v_cntr_reg(8) = '0' and v_cntr_reg(3) = '1')))) else
--              (others=>'0');
                
--  vga_blue <= h_cntr_reg(5 downto 2) when (active = '1' and ((h_cntr_reg < 512 and v_cntr_reg < 256) and  h_cntr_reg(6) = '1')) else
--              (others=>'1')          when (active = '1' and ((h_cntr_reg < 512 and not(v_cntr_reg < 256)) and not(pixel_in_box = '1'))) else 
--              (others=>'1')          when (active = '1' and ((not(h_cntr_reg < 512) and (v_cntr_reg(8) = '1' and h_cntr_reg(3) = '1')) or
--                                           (not(h_cntr_reg < 512) and (v_cntr_reg(8) = '0' and v_cntr_reg(3) = '1')))) else
--              (others=>'0');  
              
--  vga_green <= h_cntr_reg(5 downto 2) when (active = '1' and ((h_cntr_reg < 512 and v_cntr_reg < 256) and h_cntr_reg(7) = '1')) else
--              (others=>'1')           when (active = '1' and ((h_cntr_reg < 512 and not(v_cntr_reg < 256)) and not(pixel_in_box = '1'))) else 
--              (others=>'1')           when (active = '1' and ((not(h_cntr_reg < 512) and (v_cntr_reg(8) = '1' and h_cntr_reg(3) = '1')) or
--                                            (not(h_cntr_reg < 512) and (v_cntr_reg(8) = '0' and v_cntr_reg(3) = '1')))) else
--              (others=>'0');
              
 
 ------------------------------------------------------
 -------         SYNC GENERATION                 ------
 ------------------------------------------------------
 
  process (pxl_clk)
  begin
    if (rising_edge(pxl_clk)) then
      if (h_cntr_reg = (H_MAX - 1)) then
        h_cntr_reg <= (others =>'0');
      else
        h_cntr_reg <= h_cntr_reg + 1;
      end if;
    end if;
  end process;
  
  process (pxl_clk)
  begin
    if (rising_edge(pxl_clk)) then
      if ((h_cntr_reg = (H_MAX - 1)) and (v_cntr_reg = (V_MAX - 1))) then
        v_cntr_reg <= (others =>'0');
      elsif (h_cntr_reg = (H_MAX - 1)) then
        v_cntr_reg <= v_cntr_reg + 1;
      end if;
    end if;
  end process;
  
  process (pxl_clk)
  begin
    if (rising_edge(pxl_clk)) then
      if (h_cntr_reg >= (H_FP + FRAME_WIDTH - 1)) and (h_cntr_reg < (H_FP + FRAME_WIDTH + H_PW - 1)) then
        h_sync_reg <= H_POL;
      else
        h_sync_reg <= not(H_POL);
      end if;
    end if;
  end process;
  
  
  process (pxl_clk)
  begin
    if (rising_edge(pxl_clk)) then
      if (v_cntr_reg >= (V_FP + FRAME_HEIGHT - 1)) and (v_cntr_reg < (V_FP + FRAME_HEIGHT + V_PW - 1)) then
        v_sync_reg <= V_POL;
      else
        v_sync_reg <= not(V_POL);
      end if;
    end if;
  end process;
  
  
--  active <= '1' when ((h_cntr_reg < FRAME_WIDTH) and (v_cntr_reg < FRAME_HEIGHT))else
--            '0';
--active <= '1' when h_cntr_reg >= FIRST_COL and h_cntr_reg < LAST_COL and v_cntr_reg >= FIRST_LINE and v_cntr_reg < LAST_LINE else
--          '0'; 

--active <= '1' when h_cntr_reg <= FRAME_WIDTH and v_cntr_reg <= FRAME_HEIGHT else
--          '0'; 
--signal active : std_logic := '0';
  process (pxl_clk)
  begin
    if (rising_edge(pxl_clk)) then
      if(h_cntr_reg < FRAME_WIDTH and v_cntr_reg < FRAME_HEIGHT - FRAME_H_START  and v_cntr_reg >= FRAME_H_START) then
        active <='1';
      else
        active <='0';
      end if;
    end if;
  end process;
  process (pxl_clk)
  begin
    if (rising_edge(pxl_clk)) then
      v_sync_dly_reg <= v_sync_reg;
      h_sync_dly_reg <= h_sync_reg;
--      vga_red_reg <= vga_red;
--      vga_green_reg <= vga_green;
--      vga_blue_reg <= vga_blue;
    end if;
  end process;

  process (pxl_clk)
  begin
    if (rising_edge(pxl_clk)) then
	    if (h_cntr_reg < FRAME_WIDTH and v_cntr_reg < FRAME_HEIGHT - FRAME_H_START and v_cntr_reg >= FRAME_H_START) then
		  pxl_adr <= pxl_adr + 1;
		elsif ((h_cntr_reg = (H_MAX - 1)) and (v_cntr_reg = (V_MAX - 1))) then
		  pxl_adr <= (others=>'0');
		else
		  pxl_adr <= pxl_adr; 
		end if;
	end if;

--    if (rising_edge(pxl_clk)) then
--        --if (h_cntr_reg >= FIRST_COL - 1 and h_cntr_reg < LAST_COL - 1 and v_cntr_reg >= FIRST_LINE and v_cntr_reg < LAST_LINE ) then
--		if ( active = '1' ) then
--          pxl_adr <= pxl_adr + 1;
--        elsif((h_cntr_reg = (H_MAX - 2)) and (v_cntr_reg = (V_MAX - 1))) then
--          pxl_adr <= (others=>'0'); 
--        else 
--          pxl_adr <= pxl_adr; 
--        end if;
--    end if;
  end process;
  
  PXL_ADR_O <= pxl_adr;
  
  VGA_HS_O <= h_sync_dly_reg;
  VGA_VS_O <= v_sync_dly_reg;
  
  VGA_R <=PIXEL_I(7 downto 5) & "0" when active = '1' else (others=>'0');
  VGA_G <=PIXEL_I(4 downto 2) & "0" when active = '1' else (others=>'0');
  VGA_B <= PIXEL_I(1 downto 0) & "00"when active = '1' else (others=>'0');
--       /* assign VGA_R = active_s==1'b1 ? {dataout[7:5],1'b0} : 4'd0;
--   assign VGA_G = active_s==1'b1 ? {dataout[4:2],1'b0}  : 4'd0;
--   assign VGA_B = active_s==1'b1 ? {dataout[1:0],2'b00} : 4'd0;     
--   */

--  VGA_G <= vga_green_reg;
--  VGA_B <= vga_blue_reg;

end Behavioral;
