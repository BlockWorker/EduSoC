`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: University of Stuttgart, ITI
// Engineer: 
// 
// License: CERN-OHL-W-2.0
// 
// Create Date:
// Design Name: 
// Module Name: MUX_4x1_32
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module MUX_4x1_32 (
    input  [31:0] I0,
    input  [31:0] I1,
    input  [31:0] I2,
    input  [31:0] I3,
    input  [ 1:0] S,
    output [31:0] Y
);

  assign Y = S[1] ? (S[0] ? I3 : I2) : (S[0] ? I1 : I0);
endmodule
